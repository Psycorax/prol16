--------------------------------------------------------------------------------
-- Title       : 
-- Project     : 
--------------------------------------------------------------------------------
-- RevCtrl     : 
-- Authors     : 
--------------------------------------------------------------------------------
-- Description : 
--------------------------------------------------------------------------------

architecture Rtl of alu is

begin

end RTL;
