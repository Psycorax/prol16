--------------------------------------------------------------------------------
-- Title       : 
-- Project     : 
--------------------------------------------------------------------------------
-- RevCtrl     : 
-- Authors     : 
--------------------------------------------------------------------------------
-- Description : 
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- use work.Global.all;

entity DspSyncChannels is

  generic (
    
    );

  port (

    );

end DspSyncChannels;

