--------------------------------------------------------------------------------
-- Title       :
-- Project     : 
--------------------------------------------------------------------------------
-- RevCtrl     : 
-- Authors     : 
--------------------------------------------------------------------------------
-- Description : 
--------------------------------------------------------------------------------

library std;
use std.textio.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library modelsim_lib;
use modelsim_lib.util.all;

library work;
use work.prol16_pack.all;

entity tbTempl is
end tbTempl;

architecture Bhv of tbTempl is

begin

end Bhv;
